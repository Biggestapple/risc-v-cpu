library verilog;
use verilog.vl_types.all;
entity soc_ez_tb is
end soc_ez_tb;
